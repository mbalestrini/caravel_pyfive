VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pyfive_top
  CLASS BLOCK ;
  FOREIGN pyfive_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 2270.680 BY 1367.170 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 203.295 10.640 204.895 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.295 501.680 204.895 865.490 ;
    END
    PORT
      LAYER met4 ;
        RECT 203.295 1271.350 204.895 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 468.445 10.640 470.045 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 468.445 501.680 470.045 865.490 ;
    END
    PORT
      LAYER met4 ;
        RECT 468.445 1271.350 470.045 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.595 10.640 735.195 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.595 501.680 735.195 865.490 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.595 1271.350 735.195 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.745 10.640 1000.345 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.745 501.680 1000.345 865.490 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.745 1271.350 1000.345 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.895 10.640 1265.495 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.895 501.680 1265.495 865.490 ;
    END
    PORT
      LAYER met4 ;
        RECT 1263.895 1271.350 1265.495 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1529.045 10.640 1530.645 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 1529.045 501.680 1530.645 865.490 ;
    END
    PORT
      LAYER met4 ;
        RECT 1529.045 1271.350 1530.645 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1794.195 10.640 1795.795 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 1794.195 501.680 1795.795 865.490 ;
    END
    PORT
      LAYER met4 ;
        RECT 1794.195 1271.350 1795.795 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2059.345 10.640 2060.945 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 2059.345 501.680 2060.945 865.490 ;
    END
    PORT
      LAYER met4 ;
        RECT 2059.345 1271.350 2060.945 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.580 86.800 48.180 511.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.100 859.280 605.700 1278.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.580 859.280 48.180 1278.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.100 86.800 605.700 511.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1134.020 86.800 1135.620 511.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1664.860 859.280 1666.460 1278.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1134.020 859.280 1135.620 1278.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 1664.860 86.800 1666.460 511.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2222.380 86.800 2223.980 511.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2222.380 859.280 2223.980 1278.640 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 70.720 10.640 72.320 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 335.870 10.640 337.470 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 335.870 501.680 337.470 864.870 ;
    END
    PORT
      LAYER met4 ;
        RECT 335.870 1271.350 337.470 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 601.020 10.640 602.620 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 866.170 10.640 867.770 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 866.170 501.680 867.770 864.870 ;
    END
    PORT
      LAYER met4 ;
        RECT 866.170 1271.350 867.770 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1131.320 10.640 1132.920 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.470 10.640 1398.070 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.470 501.680 1398.070 864.870 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.470 1271.350 1398.070 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1661.620 10.640 1663.220 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.770 10.640 1928.370 95.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.770 501.680 1928.370 864.870 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.770 1271.350 1928.370 1354.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2191.920 10.640 2193.520 1354.800 ;
    END
  END VPWR
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 27.920 2270.680 28.520 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 864.320 2270.680 864.920 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 947.960 2270.680 948.560 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1031.600 2270.680 1032.200 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1115.240 2270.680 1115.840 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1198.880 2270.680 1199.480 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1282.520 2270.680 1283.120 ;
    END
  END io_in[15]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 111.560 2270.680 112.160 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 195.200 2270.680 195.800 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 278.840 2270.680 279.440 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 362.480 2270.680 363.080 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 446.120 2270.680 446.720 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 529.760 2270.680 530.360 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 613.400 2270.680 614.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 697.040 2270.680 697.640 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 780.680 2270.680 781.280 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 55.800 2270.680 56.400 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 892.200 2270.680 892.800 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 975.840 2270.680 976.440 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1059.480 2270.680 1060.080 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1143.120 2270.680 1143.720 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1226.760 2270.680 1227.360 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1310.400 2270.680 1311.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 139.440 2270.680 140.040 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 223.080 2270.680 223.680 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 306.720 2270.680 307.320 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 390.360 2270.680 390.960 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 474.000 2270.680 474.600 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 557.640 2270.680 558.240 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 641.280 2270.680 641.880 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 724.920 2270.680 725.520 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 808.560 2270.680 809.160 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 83.680 2270.680 84.280 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 920.080 2270.680 920.680 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1003.720 2270.680 1004.320 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1087.360 2270.680 1087.960 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1171.000 2270.680 1171.600 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1254.640 2270.680 1255.240 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 1338.280 2270.680 1338.880 ;
    END
  END io_out[15]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 167.320 2270.680 167.920 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 250.960 2270.680 251.560 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 334.600 2270.680 335.200 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 418.240 2270.680 418.840 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 501.880 2270.680 502.480 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 585.520 2270.680 586.120 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 669.160 2270.680 669.760 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 752.800 2270.680 753.400 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2266.680 836.440 2270.680 837.040 ;
    END
  END io_out[9]
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.550 1363.170 1702.830 1367.170 ;
    END
  END one
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.760 4.000 530.360 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 566.480 4.000 567.080 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.200 4.000 603.800 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 713.360 4.000 713.960 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.080 4.000 750.680 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.800 4.000 787.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 823.520 4.000 824.120 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.240 4.000 860.840 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.960 4.000 897.560 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.680 4.000 934.280 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 970.400 4.000 971.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.120 4.000 1007.720 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1043.840 4.000 1044.440 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1080.560 4.000 1081.160 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1117.280 4.000 1117.880 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1154.000 4.000 1154.600 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.720 4.000 1191.320 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1264.160 4.000 1264.760 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1300.880 4.000 1301.480 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.600 4.000 420.200 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 456.320 4.000 456.920 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.000 4.000 542.600 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 725.600 4.000 726.200 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 762.320 4.000 762.920 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.760 4.000 836.360 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 872.480 4.000 873.080 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.200 4.000 909.800 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.920 4.000 946.520 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 982.640 4.000 983.240 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1019.360 4.000 1019.960 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.080 4.000 1056.680 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1092.800 4.000 1093.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1129.520 4.000 1130.120 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1166.240 4.000 1166.840 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1202.960 4.000 1203.560 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1239.680 4.000 1240.280 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1276.400 4.000 1277.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1313.120 4.000 1313.720 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.720 4.000 273.320 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.280 4.000 505.880 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.680 4.000 628.280 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 664.400 4.000 665.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.120 4.000 701.720 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 774.560 4.000 775.160 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.280 4.000 811.880 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.000 4.000 848.600 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.720 4.000 885.320 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.160 4.000 958.760 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.880 4.000 995.480 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1031.600 4.000 1032.200 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1068.320 4.000 1068.920 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1105.040 4.000 1105.640 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.760 4.000 1142.360 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1178.480 4.000 1179.080 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1215.200 4.000 1215.800 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1251.920 4.000 1252.520 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1288.640 4.000 1289.240 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1325.360 4.000 1325.960 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.960 4.000 285.560 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.920 4.000 334.520 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 517.520 4.000 518.120 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.320 4.000 150.920 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END wbs_we_i
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 1363.170 567.550 1367.170 ;
    END
  END zero
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2265.040 1354.645 ;
      LAYER met1 ;
        RECT 5.520 10.640 2265.040 1354.800 ;
      LAYER met2 ;
        RECT 7.000 1362.890 566.990 1363.810 ;
        RECT 567.830 1362.890 1702.270 1363.810 ;
        RECT 1703.110 1362.890 2262.650 1363.810 ;
        RECT 7.000 10.695 2262.650 1362.890 ;
      LAYER met3 ;
        RECT 4.000 1339.280 2266.680 1354.725 ;
        RECT 4.000 1337.880 2266.280 1339.280 ;
        RECT 4.000 1326.360 2266.680 1337.880 ;
        RECT 4.400 1324.960 2266.680 1326.360 ;
        RECT 4.000 1314.120 2266.680 1324.960 ;
        RECT 4.400 1312.720 2266.680 1314.120 ;
        RECT 4.000 1311.400 2266.680 1312.720 ;
        RECT 4.000 1310.000 2266.280 1311.400 ;
        RECT 4.000 1301.880 2266.680 1310.000 ;
        RECT 4.400 1300.480 2266.680 1301.880 ;
        RECT 4.000 1289.640 2266.680 1300.480 ;
        RECT 4.400 1288.240 2266.680 1289.640 ;
        RECT 4.000 1283.520 2266.680 1288.240 ;
        RECT 4.000 1282.120 2266.280 1283.520 ;
        RECT 4.000 1277.400 2266.680 1282.120 ;
        RECT 4.400 1276.000 2266.680 1277.400 ;
        RECT 4.000 1265.160 2266.680 1276.000 ;
        RECT 4.400 1263.760 2266.680 1265.160 ;
        RECT 4.000 1255.640 2266.680 1263.760 ;
        RECT 4.000 1254.240 2266.280 1255.640 ;
        RECT 4.000 1252.920 2266.680 1254.240 ;
        RECT 4.400 1251.520 2266.680 1252.920 ;
        RECT 4.000 1240.680 2266.680 1251.520 ;
        RECT 4.400 1239.280 2266.680 1240.680 ;
        RECT 4.000 1228.440 2266.680 1239.280 ;
        RECT 4.400 1227.760 2266.680 1228.440 ;
        RECT 4.400 1227.040 2266.280 1227.760 ;
        RECT 4.000 1226.360 2266.280 1227.040 ;
        RECT 4.000 1216.200 2266.680 1226.360 ;
        RECT 4.400 1214.800 2266.680 1216.200 ;
        RECT 4.000 1203.960 2266.680 1214.800 ;
        RECT 4.400 1202.560 2266.680 1203.960 ;
        RECT 4.000 1199.880 2266.680 1202.560 ;
        RECT 4.000 1198.480 2266.280 1199.880 ;
        RECT 4.000 1191.720 2266.680 1198.480 ;
        RECT 4.400 1190.320 2266.680 1191.720 ;
        RECT 4.000 1179.480 2266.680 1190.320 ;
        RECT 4.400 1178.080 2266.680 1179.480 ;
        RECT 4.000 1172.000 2266.680 1178.080 ;
        RECT 4.000 1170.600 2266.280 1172.000 ;
        RECT 4.000 1167.240 2266.680 1170.600 ;
        RECT 4.400 1165.840 2266.680 1167.240 ;
        RECT 4.000 1155.000 2266.680 1165.840 ;
        RECT 4.400 1153.600 2266.680 1155.000 ;
        RECT 4.000 1144.120 2266.680 1153.600 ;
        RECT 4.000 1142.760 2266.280 1144.120 ;
        RECT 4.400 1142.720 2266.280 1142.760 ;
        RECT 4.400 1141.360 2266.680 1142.720 ;
        RECT 4.000 1130.520 2266.680 1141.360 ;
        RECT 4.400 1129.120 2266.680 1130.520 ;
        RECT 4.000 1118.280 2266.680 1129.120 ;
        RECT 4.400 1116.880 2266.680 1118.280 ;
        RECT 4.000 1116.240 2266.680 1116.880 ;
        RECT 4.000 1114.840 2266.280 1116.240 ;
        RECT 4.000 1106.040 2266.680 1114.840 ;
        RECT 4.400 1104.640 2266.680 1106.040 ;
        RECT 4.000 1093.800 2266.680 1104.640 ;
        RECT 4.400 1092.400 2266.680 1093.800 ;
        RECT 4.000 1088.360 2266.680 1092.400 ;
        RECT 4.000 1086.960 2266.280 1088.360 ;
        RECT 4.000 1081.560 2266.680 1086.960 ;
        RECT 4.400 1080.160 2266.680 1081.560 ;
        RECT 4.000 1069.320 2266.680 1080.160 ;
        RECT 4.400 1067.920 2266.680 1069.320 ;
        RECT 4.000 1060.480 2266.680 1067.920 ;
        RECT 4.000 1059.080 2266.280 1060.480 ;
        RECT 4.000 1057.080 2266.680 1059.080 ;
        RECT 4.400 1055.680 2266.680 1057.080 ;
        RECT 4.000 1044.840 2266.680 1055.680 ;
        RECT 4.400 1043.440 2266.680 1044.840 ;
        RECT 4.000 1032.600 2266.680 1043.440 ;
        RECT 4.400 1031.200 2266.280 1032.600 ;
        RECT 4.000 1020.360 2266.680 1031.200 ;
        RECT 4.400 1018.960 2266.680 1020.360 ;
        RECT 4.000 1008.120 2266.680 1018.960 ;
        RECT 4.400 1006.720 2266.680 1008.120 ;
        RECT 4.000 1004.720 2266.680 1006.720 ;
        RECT 4.000 1003.320 2266.280 1004.720 ;
        RECT 4.000 995.880 2266.680 1003.320 ;
        RECT 4.400 994.480 2266.680 995.880 ;
        RECT 4.000 983.640 2266.680 994.480 ;
        RECT 4.400 982.240 2266.680 983.640 ;
        RECT 4.000 976.840 2266.680 982.240 ;
        RECT 4.000 975.440 2266.280 976.840 ;
        RECT 4.000 971.400 2266.680 975.440 ;
        RECT 4.400 970.000 2266.680 971.400 ;
        RECT 4.000 959.160 2266.680 970.000 ;
        RECT 4.400 957.760 2266.680 959.160 ;
        RECT 4.000 948.960 2266.680 957.760 ;
        RECT 4.000 947.560 2266.280 948.960 ;
        RECT 4.000 946.920 2266.680 947.560 ;
        RECT 4.400 945.520 2266.680 946.920 ;
        RECT 4.000 934.680 2266.680 945.520 ;
        RECT 4.400 933.280 2266.680 934.680 ;
        RECT 4.000 922.440 2266.680 933.280 ;
        RECT 4.400 921.080 2266.680 922.440 ;
        RECT 4.400 921.040 2266.280 921.080 ;
        RECT 4.000 919.680 2266.280 921.040 ;
        RECT 4.000 910.200 2266.680 919.680 ;
        RECT 4.400 908.800 2266.680 910.200 ;
        RECT 4.000 897.960 2266.680 908.800 ;
        RECT 4.400 896.560 2266.680 897.960 ;
        RECT 4.000 893.200 2266.680 896.560 ;
        RECT 4.000 891.800 2266.280 893.200 ;
        RECT 4.000 885.720 2266.680 891.800 ;
        RECT 4.400 884.320 2266.680 885.720 ;
        RECT 4.000 873.480 2266.680 884.320 ;
        RECT 4.400 872.080 2266.680 873.480 ;
        RECT 4.000 865.320 2266.680 872.080 ;
        RECT 4.000 863.920 2266.280 865.320 ;
        RECT 4.000 861.240 2266.680 863.920 ;
        RECT 4.400 859.840 2266.680 861.240 ;
        RECT 4.000 849.000 2266.680 859.840 ;
        RECT 4.400 847.600 2266.680 849.000 ;
        RECT 4.000 837.440 2266.680 847.600 ;
        RECT 4.000 836.760 2266.280 837.440 ;
        RECT 4.400 836.040 2266.280 836.760 ;
        RECT 4.400 835.360 2266.680 836.040 ;
        RECT 4.000 824.520 2266.680 835.360 ;
        RECT 4.400 823.120 2266.680 824.520 ;
        RECT 4.000 812.280 2266.680 823.120 ;
        RECT 4.400 810.880 2266.680 812.280 ;
        RECT 4.000 809.560 2266.680 810.880 ;
        RECT 4.000 808.160 2266.280 809.560 ;
        RECT 4.000 800.040 2266.680 808.160 ;
        RECT 4.400 798.640 2266.680 800.040 ;
        RECT 4.000 787.800 2266.680 798.640 ;
        RECT 4.400 786.400 2266.680 787.800 ;
        RECT 4.000 781.680 2266.680 786.400 ;
        RECT 4.000 780.280 2266.280 781.680 ;
        RECT 4.000 775.560 2266.680 780.280 ;
        RECT 4.400 774.160 2266.680 775.560 ;
        RECT 4.000 763.320 2266.680 774.160 ;
        RECT 4.400 761.920 2266.680 763.320 ;
        RECT 4.000 753.800 2266.680 761.920 ;
        RECT 4.000 752.400 2266.280 753.800 ;
        RECT 4.000 751.080 2266.680 752.400 ;
        RECT 4.400 749.680 2266.680 751.080 ;
        RECT 4.000 738.840 2266.680 749.680 ;
        RECT 4.400 737.440 2266.680 738.840 ;
        RECT 4.000 726.600 2266.680 737.440 ;
        RECT 4.400 725.920 2266.680 726.600 ;
        RECT 4.400 725.200 2266.280 725.920 ;
        RECT 4.000 724.520 2266.280 725.200 ;
        RECT 4.000 714.360 2266.680 724.520 ;
        RECT 4.400 712.960 2266.680 714.360 ;
        RECT 4.000 702.120 2266.680 712.960 ;
        RECT 4.400 700.720 2266.680 702.120 ;
        RECT 4.000 698.040 2266.680 700.720 ;
        RECT 4.000 696.640 2266.280 698.040 ;
        RECT 4.000 689.880 2266.680 696.640 ;
        RECT 4.400 688.480 2266.680 689.880 ;
        RECT 4.000 677.640 2266.680 688.480 ;
        RECT 4.400 676.240 2266.680 677.640 ;
        RECT 4.000 670.160 2266.680 676.240 ;
        RECT 4.000 668.760 2266.280 670.160 ;
        RECT 4.000 665.400 2266.680 668.760 ;
        RECT 4.400 664.000 2266.680 665.400 ;
        RECT 4.000 653.160 2266.680 664.000 ;
        RECT 4.400 651.760 2266.680 653.160 ;
        RECT 4.000 642.280 2266.680 651.760 ;
        RECT 4.000 640.920 2266.280 642.280 ;
        RECT 4.400 640.880 2266.280 640.920 ;
        RECT 4.400 639.520 2266.680 640.880 ;
        RECT 4.000 628.680 2266.680 639.520 ;
        RECT 4.400 627.280 2266.680 628.680 ;
        RECT 4.000 616.440 2266.680 627.280 ;
        RECT 4.400 615.040 2266.680 616.440 ;
        RECT 4.000 614.400 2266.680 615.040 ;
        RECT 4.000 613.000 2266.280 614.400 ;
        RECT 4.000 604.200 2266.680 613.000 ;
        RECT 4.400 602.800 2266.680 604.200 ;
        RECT 4.000 591.960 2266.680 602.800 ;
        RECT 4.400 590.560 2266.680 591.960 ;
        RECT 4.000 586.520 2266.680 590.560 ;
        RECT 4.000 585.120 2266.280 586.520 ;
        RECT 4.000 579.720 2266.680 585.120 ;
        RECT 4.400 578.320 2266.680 579.720 ;
        RECT 4.000 567.480 2266.680 578.320 ;
        RECT 4.400 566.080 2266.680 567.480 ;
        RECT 4.000 558.640 2266.680 566.080 ;
        RECT 4.000 557.240 2266.280 558.640 ;
        RECT 4.000 555.240 2266.680 557.240 ;
        RECT 4.400 553.840 2266.680 555.240 ;
        RECT 4.000 543.000 2266.680 553.840 ;
        RECT 4.400 541.600 2266.680 543.000 ;
        RECT 4.000 530.760 2266.680 541.600 ;
        RECT 4.400 529.360 2266.280 530.760 ;
        RECT 4.000 518.520 2266.680 529.360 ;
        RECT 4.400 517.120 2266.680 518.520 ;
        RECT 4.000 506.280 2266.680 517.120 ;
        RECT 4.400 504.880 2266.680 506.280 ;
        RECT 4.000 502.880 2266.680 504.880 ;
        RECT 4.000 501.480 2266.280 502.880 ;
        RECT 4.000 494.040 2266.680 501.480 ;
        RECT 4.400 492.640 2266.680 494.040 ;
        RECT 4.000 481.800 2266.680 492.640 ;
        RECT 4.400 480.400 2266.680 481.800 ;
        RECT 4.000 475.000 2266.680 480.400 ;
        RECT 4.000 473.600 2266.280 475.000 ;
        RECT 4.000 469.560 2266.680 473.600 ;
        RECT 4.400 468.160 2266.680 469.560 ;
        RECT 4.000 457.320 2266.680 468.160 ;
        RECT 4.400 455.920 2266.680 457.320 ;
        RECT 4.000 447.120 2266.680 455.920 ;
        RECT 4.000 445.720 2266.280 447.120 ;
        RECT 4.000 445.080 2266.680 445.720 ;
        RECT 4.400 443.680 2266.680 445.080 ;
        RECT 4.000 432.840 2266.680 443.680 ;
        RECT 4.400 431.440 2266.680 432.840 ;
        RECT 4.000 420.600 2266.680 431.440 ;
        RECT 4.400 419.240 2266.680 420.600 ;
        RECT 4.400 419.200 2266.280 419.240 ;
        RECT 4.000 417.840 2266.280 419.200 ;
        RECT 4.000 408.360 2266.680 417.840 ;
        RECT 4.400 406.960 2266.680 408.360 ;
        RECT 4.000 396.120 2266.680 406.960 ;
        RECT 4.400 394.720 2266.680 396.120 ;
        RECT 4.000 391.360 2266.680 394.720 ;
        RECT 4.000 389.960 2266.280 391.360 ;
        RECT 4.000 383.880 2266.680 389.960 ;
        RECT 4.400 382.480 2266.680 383.880 ;
        RECT 4.000 371.640 2266.680 382.480 ;
        RECT 4.400 370.240 2266.680 371.640 ;
        RECT 4.000 363.480 2266.680 370.240 ;
        RECT 4.000 362.080 2266.280 363.480 ;
        RECT 4.000 359.400 2266.680 362.080 ;
        RECT 4.400 358.000 2266.680 359.400 ;
        RECT 4.000 347.160 2266.680 358.000 ;
        RECT 4.400 345.760 2266.680 347.160 ;
        RECT 4.000 335.600 2266.680 345.760 ;
        RECT 4.000 334.920 2266.280 335.600 ;
        RECT 4.400 334.200 2266.280 334.920 ;
        RECT 4.400 333.520 2266.680 334.200 ;
        RECT 4.000 322.680 2266.680 333.520 ;
        RECT 4.400 321.280 2266.680 322.680 ;
        RECT 4.000 310.440 2266.680 321.280 ;
        RECT 4.400 309.040 2266.680 310.440 ;
        RECT 4.000 307.720 2266.680 309.040 ;
        RECT 4.000 306.320 2266.280 307.720 ;
        RECT 4.000 298.200 2266.680 306.320 ;
        RECT 4.400 296.800 2266.680 298.200 ;
        RECT 4.000 285.960 2266.680 296.800 ;
        RECT 4.400 284.560 2266.680 285.960 ;
        RECT 4.000 279.840 2266.680 284.560 ;
        RECT 4.000 278.440 2266.280 279.840 ;
        RECT 4.000 273.720 2266.680 278.440 ;
        RECT 4.400 272.320 2266.680 273.720 ;
        RECT 4.000 261.480 2266.680 272.320 ;
        RECT 4.400 260.080 2266.680 261.480 ;
        RECT 4.000 251.960 2266.680 260.080 ;
        RECT 4.000 250.560 2266.280 251.960 ;
        RECT 4.000 249.240 2266.680 250.560 ;
        RECT 4.400 247.840 2266.680 249.240 ;
        RECT 4.000 237.000 2266.680 247.840 ;
        RECT 4.400 235.600 2266.680 237.000 ;
        RECT 4.000 224.760 2266.680 235.600 ;
        RECT 4.400 224.080 2266.680 224.760 ;
        RECT 4.400 223.360 2266.280 224.080 ;
        RECT 4.000 222.680 2266.280 223.360 ;
        RECT 4.000 212.520 2266.680 222.680 ;
        RECT 4.400 211.120 2266.680 212.520 ;
        RECT 4.000 200.280 2266.680 211.120 ;
        RECT 4.400 198.880 2266.680 200.280 ;
        RECT 4.000 196.200 2266.680 198.880 ;
        RECT 4.000 194.800 2266.280 196.200 ;
        RECT 4.000 188.040 2266.680 194.800 ;
        RECT 4.400 186.640 2266.680 188.040 ;
        RECT 4.000 175.800 2266.680 186.640 ;
        RECT 4.400 174.400 2266.680 175.800 ;
        RECT 4.000 168.320 2266.680 174.400 ;
        RECT 4.000 166.920 2266.280 168.320 ;
        RECT 4.000 163.560 2266.680 166.920 ;
        RECT 4.400 162.160 2266.680 163.560 ;
        RECT 4.000 151.320 2266.680 162.160 ;
        RECT 4.400 149.920 2266.680 151.320 ;
        RECT 4.000 140.440 2266.680 149.920 ;
        RECT 4.000 139.080 2266.280 140.440 ;
        RECT 4.400 139.040 2266.280 139.080 ;
        RECT 4.400 137.680 2266.680 139.040 ;
        RECT 4.000 126.840 2266.680 137.680 ;
        RECT 4.400 125.440 2266.680 126.840 ;
        RECT 4.000 114.600 2266.680 125.440 ;
        RECT 4.400 113.200 2266.680 114.600 ;
        RECT 4.000 112.560 2266.680 113.200 ;
        RECT 4.000 111.160 2266.280 112.560 ;
        RECT 4.000 102.360 2266.680 111.160 ;
        RECT 4.400 100.960 2266.680 102.360 ;
        RECT 4.000 90.120 2266.680 100.960 ;
        RECT 4.400 88.720 2266.680 90.120 ;
        RECT 4.000 84.680 2266.680 88.720 ;
        RECT 4.000 83.280 2266.280 84.680 ;
        RECT 4.000 77.880 2266.680 83.280 ;
        RECT 4.400 76.480 2266.680 77.880 ;
        RECT 4.000 65.640 2266.680 76.480 ;
        RECT 4.400 64.240 2266.680 65.640 ;
        RECT 4.000 56.800 2266.680 64.240 ;
        RECT 4.000 55.400 2266.280 56.800 ;
        RECT 4.000 53.400 2266.680 55.400 ;
        RECT 4.400 52.000 2266.680 53.400 ;
        RECT 4.000 41.160 2266.680 52.000 ;
        RECT 4.400 39.760 2266.680 41.160 ;
        RECT 4.000 28.920 2266.680 39.760 ;
        RECT 4.000 27.520 2266.280 28.920 ;
        RECT 4.000 10.715 2266.680 27.520 ;
      LAYER met4 ;
        RECT 78.495 1270.950 202.895 1285.705 ;
        RECT 205.295 1270.950 335.470 1285.705 ;
        RECT 337.870 1270.950 468.045 1285.705 ;
        RECT 470.445 1270.950 600.620 1285.705 ;
        RECT 78.495 865.890 600.620 1270.950 ;
        RECT 78.495 501.280 202.895 865.890 ;
        RECT 205.295 865.270 468.045 865.890 ;
        RECT 205.295 501.280 335.470 865.270 ;
        RECT 337.870 501.280 468.045 865.270 ;
        RECT 470.445 501.280 600.620 865.890 ;
        RECT 78.495 96.220 600.620 501.280 ;
        RECT 78.495 39.615 202.895 96.220 ;
        RECT 205.295 39.615 335.470 96.220 ;
        RECT 337.870 39.615 468.045 96.220 ;
        RECT 470.445 39.615 600.620 96.220 ;
        RECT 603.020 1279.040 733.195 1285.705 ;
        RECT 603.020 858.880 603.700 1279.040 ;
        RECT 606.100 1270.950 733.195 1279.040 ;
        RECT 735.595 1270.950 865.770 1285.705 ;
        RECT 868.170 1270.950 998.345 1285.705 ;
        RECT 1000.745 1270.950 1130.920 1285.705 ;
        RECT 606.100 865.890 1130.920 1270.950 ;
        RECT 606.100 858.880 733.195 865.890 ;
        RECT 603.020 512.000 733.195 858.880 ;
        RECT 603.020 86.400 603.700 512.000 ;
        RECT 606.100 501.280 733.195 512.000 ;
        RECT 735.595 865.270 998.345 865.890 ;
        RECT 735.595 501.280 865.770 865.270 ;
        RECT 868.170 501.280 998.345 865.270 ;
        RECT 1000.745 501.280 1130.920 865.890 ;
        RECT 606.100 96.220 1130.920 501.280 ;
        RECT 606.100 86.400 733.195 96.220 ;
        RECT 603.020 39.615 733.195 86.400 ;
        RECT 735.595 39.615 865.770 96.220 ;
        RECT 868.170 39.615 998.345 96.220 ;
        RECT 1000.745 39.615 1130.920 96.220 ;
        RECT 1133.320 1279.040 1263.495 1285.705 ;
        RECT 1133.320 858.880 1133.620 1279.040 ;
        RECT 1136.020 1270.950 1263.495 1279.040 ;
        RECT 1265.895 1270.950 1396.070 1285.705 ;
        RECT 1398.470 1270.950 1528.645 1285.705 ;
        RECT 1531.045 1270.950 1661.220 1285.705 ;
        RECT 1136.020 865.890 1661.220 1270.950 ;
        RECT 1136.020 858.880 1263.495 865.890 ;
        RECT 1133.320 512.000 1263.495 858.880 ;
        RECT 1133.320 86.400 1133.620 512.000 ;
        RECT 1136.020 501.280 1263.495 512.000 ;
        RECT 1265.895 865.270 1528.645 865.890 ;
        RECT 1265.895 501.280 1396.070 865.270 ;
        RECT 1398.470 501.280 1528.645 865.270 ;
        RECT 1531.045 501.280 1661.220 865.890 ;
        RECT 1136.020 96.220 1661.220 501.280 ;
        RECT 1136.020 86.400 1263.495 96.220 ;
        RECT 1133.320 39.615 1263.495 86.400 ;
        RECT 1265.895 39.615 1396.070 96.220 ;
        RECT 1398.470 39.615 1528.645 96.220 ;
        RECT 1531.045 39.615 1661.220 96.220 ;
        RECT 1663.620 1279.040 1793.795 1285.705 ;
        RECT 1663.620 858.880 1664.460 1279.040 ;
        RECT 1666.860 1270.950 1793.795 1279.040 ;
        RECT 1796.195 1270.950 1926.370 1285.705 ;
        RECT 1928.770 1270.950 2058.945 1285.705 ;
        RECT 2061.345 1270.950 2187.465 1285.705 ;
        RECT 1666.860 865.890 2187.465 1270.950 ;
        RECT 1666.860 858.880 1793.795 865.890 ;
        RECT 1663.620 512.000 1793.795 858.880 ;
        RECT 1663.620 86.400 1664.460 512.000 ;
        RECT 1666.860 501.280 1793.795 512.000 ;
        RECT 1796.195 865.270 2058.945 865.890 ;
        RECT 1796.195 501.280 1926.370 865.270 ;
        RECT 1928.770 501.280 2058.945 865.270 ;
        RECT 2061.345 501.280 2187.465 865.890 ;
        RECT 1666.860 96.220 2187.465 501.280 ;
        RECT 1666.860 86.400 1793.795 96.220 ;
        RECT 1663.620 39.615 1793.795 86.400 ;
        RECT 1796.195 39.615 1926.370 96.220 ;
        RECT 1928.770 39.615 2058.945 96.220 ;
        RECT 2061.345 39.615 2187.465 96.220 ;
  END
END pyfive_top
END LIBRARY

