magic
tech sky130A
magscale 1 2
timestamp 1672422764
<< obsli1 >>
rect 1104 2159 453008 270929
<< obsm1 >>
rect 1104 2128 453008 270960
<< metal2 >>
rect 113454 272634 113510 273434
rect 340510 272634 340566 273434
<< obsm2 >>
rect 1400 272578 113398 272762
rect 113566 272578 340454 272762
rect 340622 272578 452530 272762
rect 1400 2139 452530 272578
<< metal3 >>
rect 453336 267656 454136 267776
rect 0 265072 800 265192
rect 0 262624 800 262744
rect 453336 262080 454136 262200
rect 0 260176 800 260296
rect 0 257728 800 257848
rect 453336 256504 454136 256624
rect 0 255280 800 255400
rect 0 252832 800 252952
rect 453336 250928 454136 251048
rect 0 250384 800 250504
rect 0 247936 800 248056
rect 0 245488 800 245608
rect 453336 245352 454136 245472
rect 0 243040 800 243160
rect 0 240592 800 240712
rect 453336 239776 454136 239896
rect 0 238144 800 238264
rect 0 235696 800 235816
rect 453336 234200 454136 234320
rect 0 233248 800 233368
rect 0 230800 800 230920
rect 453336 228624 454136 228744
rect 0 228352 800 228472
rect 0 225904 800 226024
rect 0 223456 800 223576
rect 453336 223048 454136 223168
rect 0 221008 800 221128
rect 0 218560 800 218680
rect 453336 217472 454136 217592
rect 0 216112 800 216232
rect 0 213664 800 213784
rect 453336 211896 454136 212016
rect 0 211216 800 211336
rect 0 208768 800 208888
rect 0 206320 800 206440
rect 453336 206320 454136 206440
rect 0 203872 800 203992
rect 0 201424 800 201544
rect 453336 200744 454136 200864
rect 0 198976 800 199096
rect 0 196528 800 196648
rect 453336 195168 454136 195288
rect 0 194080 800 194200
rect 0 191632 800 191752
rect 453336 189592 454136 189712
rect 0 189184 800 189304
rect 0 186736 800 186856
rect 0 184288 800 184408
rect 453336 184016 454136 184136
rect 0 181840 800 181960
rect 0 179392 800 179512
rect 453336 178440 454136 178560
rect 0 176944 800 177064
rect 0 174496 800 174616
rect 453336 172864 454136 172984
rect 0 172048 800 172168
rect 0 169600 800 169720
rect 0 167152 800 167272
rect 453336 167288 454136 167408
rect 0 164704 800 164824
rect 0 162256 800 162376
rect 453336 161712 454136 161832
rect 0 159808 800 159928
rect 0 157360 800 157480
rect 453336 156136 454136 156256
rect 0 154912 800 155032
rect 0 152464 800 152584
rect 453336 150560 454136 150680
rect 0 150016 800 150136
rect 0 147568 800 147688
rect 0 145120 800 145240
rect 453336 144984 454136 145104
rect 0 142672 800 142792
rect 0 140224 800 140344
rect 453336 139408 454136 139528
rect 0 137776 800 137896
rect 0 135328 800 135448
rect 453336 133832 454136 133952
rect 0 132880 800 133000
rect 0 130432 800 130552
rect 453336 128256 454136 128376
rect 0 127984 800 128104
rect 0 125536 800 125656
rect 0 123088 800 123208
rect 453336 122680 454136 122800
rect 0 120640 800 120760
rect 0 118192 800 118312
rect 453336 117104 454136 117224
rect 0 115744 800 115864
rect 0 113296 800 113416
rect 453336 111528 454136 111648
rect 0 110848 800 110968
rect 0 108400 800 108520
rect 0 105952 800 106072
rect 453336 105952 454136 106072
rect 0 103504 800 103624
rect 0 101056 800 101176
rect 453336 100376 454136 100496
rect 0 98608 800 98728
rect 0 96160 800 96280
rect 453336 94800 454136 94920
rect 0 93712 800 93832
rect 0 91264 800 91384
rect 453336 89224 454136 89344
rect 0 88816 800 88936
rect 0 86368 800 86488
rect 0 83920 800 84040
rect 453336 83648 454136 83768
rect 0 81472 800 81592
rect 0 79024 800 79144
rect 453336 78072 454136 78192
rect 0 76576 800 76696
rect 0 74128 800 74248
rect 453336 72496 454136 72616
rect 0 71680 800 71800
rect 0 69232 800 69352
rect 0 66784 800 66904
rect 453336 66920 454136 67040
rect 0 64336 800 64456
rect 0 61888 800 62008
rect 453336 61344 454136 61464
rect 0 59440 800 59560
rect 0 56992 800 57112
rect 453336 55768 454136 55888
rect 0 54544 800 54664
rect 0 52096 800 52216
rect 453336 50192 454136 50312
rect 0 49648 800 49768
rect 0 47200 800 47320
rect 0 44752 800 44872
rect 453336 44616 454136 44736
rect 0 42304 800 42424
rect 0 39856 800 39976
rect 453336 39040 454136 39160
rect 0 37408 800 37528
rect 0 34960 800 35080
rect 453336 33464 454136 33584
rect 0 32512 800 32632
rect 0 30064 800 30184
rect 453336 27888 454136 28008
rect 0 27616 800 27736
rect 0 25168 800 25288
rect 0 22720 800 22840
rect 453336 22312 454136 22432
rect 0 20272 800 20392
rect 0 17824 800 17944
rect 453336 16736 454136 16856
rect 0 15376 800 15496
rect 0 12928 800 13048
rect 453336 11160 454136 11280
rect 0 10480 800 10600
rect 0 8032 800 8152
rect 453336 5584 454136 5704
<< obsm3 >>
rect 800 267856 453336 270945
rect 800 267576 453256 267856
rect 800 265272 453336 267576
rect 880 264992 453336 265272
rect 800 262824 453336 264992
rect 880 262544 453336 262824
rect 800 262280 453336 262544
rect 800 262000 453256 262280
rect 800 260376 453336 262000
rect 880 260096 453336 260376
rect 800 257928 453336 260096
rect 880 257648 453336 257928
rect 800 256704 453336 257648
rect 800 256424 453256 256704
rect 800 255480 453336 256424
rect 880 255200 453336 255480
rect 800 253032 453336 255200
rect 880 252752 453336 253032
rect 800 251128 453336 252752
rect 800 250848 453256 251128
rect 800 250584 453336 250848
rect 880 250304 453336 250584
rect 800 248136 453336 250304
rect 880 247856 453336 248136
rect 800 245688 453336 247856
rect 880 245552 453336 245688
rect 880 245408 453256 245552
rect 800 245272 453256 245408
rect 800 243240 453336 245272
rect 880 242960 453336 243240
rect 800 240792 453336 242960
rect 880 240512 453336 240792
rect 800 239976 453336 240512
rect 800 239696 453256 239976
rect 800 238344 453336 239696
rect 880 238064 453336 238344
rect 800 235896 453336 238064
rect 880 235616 453336 235896
rect 800 234400 453336 235616
rect 800 234120 453256 234400
rect 800 233448 453336 234120
rect 880 233168 453336 233448
rect 800 231000 453336 233168
rect 880 230720 453336 231000
rect 800 228824 453336 230720
rect 800 228552 453256 228824
rect 880 228544 453256 228552
rect 880 228272 453336 228544
rect 800 226104 453336 228272
rect 880 225824 453336 226104
rect 800 223656 453336 225824
rect 880 223376 453336 223656
rect 800 223248 453336 223376
rect 800 222968 453256 223248
rect 800 221208 453336 222968
rect 880 220928 453336 221208
rect 800 218760 453336 220928
rect 880 218480 453336 218760
rect 800 217672 453336 218480
rect 800 217392 453256 217672
rect 800 216312 453336 217392
rect 880 216032 453336 216312
rect 800 213864 453336 216032
rect 880 213584 453336 213864
rect 800 212096 453336 213584
rect 800 211816 453256 212096
rect 800 211416 453336 211816
rect 880 211136 453336 211416
rect 800 208968 453336 211136
rect 880 208688 453336 208968
rect 800 206520 453336 208688
rect 880 206240 453256 206520
rect 800 204072 453336 206240
rect 880 203792 453336 204072
rect 800 201624 453336 203792
rect 880 201344 453336 201624
rect 800 200944 453336 201344
rect 800 200664 453256 200944
rect 800 199176 453336 200664
rect 880 198896 453336 199176
rect 800 196728 453336 198896
rect 880 196448 453336 196728
rect 800 195368 453336 196448
rect 800 195088 453256 195368
rect 800 194280 453336 195088
rect 880 194000 453336 194280
rect 800 191832 453336 194000
rect 880 191552 453336 191832
rect 800 189792 453336 191552
rect 800 189512 453256 189792
rect 800 189384 453336 189512
rect 880 189104 453336 189384
rect 800 186936 453336 189104
rect 880 186656 453336 186936
rect 800 184488 453336 186656
rect 880 184216 453336 184488
rect 880 184208 453256 184216
rect 800 183936 453256 184208
rect 800 182040 453336 183936
rect 880 181760 453336 182040
rect 800 179592 453336 181760
rect 880 179312 453336 179592
rect 800 178640 453336 179312
rect 800 178360 453256 178640
rect 800 177144 453336 178360
rect 880 176864 453336 177144
rect 800 174696 453336 176864
rect 880 174416 453336 174696
rect 800 173064 453336 174416
rect 800 172784 453256 173064
rect 800 172248 453336 172784
rect 880 171968 453336 172248
rect 800 169800 453336 171968
rect 880 169520 453336 169800
rect 800 167488 453336 169520
rect 800 167352 453256 167488
rect 880 167208 453256 167352
rect 880 167072 453336 167208
rect 800 164904 453336 167072
rect 880 164624 453336 164904
rect 800 162456 453336 164624
rect 880 162176 453336 162456
rect 800 161912 453336 162176
rect 800 161632 453256 161912
rect 800 160008 453336 161632
rect 880 159728 453336 160008
rect 800 157560 453336 159728
rect 880 157280 453336 157560
rect 800 156336 453336 157280
rect 800 156056 453256 156336
rect 800 155112 453336 156056
rect 880 154832 453336 155112
rect 800 152664 453336 154832
rect 880 152384 453336 152664
rect 800 150760 453336 152384
rect 800 150480 453256 150760
rect 800 150216 453336 150480
rect 880 149936 453336 150216
rect 800 147768 453336 149936
rect 880 147488 453336 147768
rect 800 145320 453336 147488
rect 880 145184 453336 145320
rect 880 145040 453256 145184
rect 800 144904 453256 145040
rect 800 142872 453336 144904
rect 880 142592 453336 142872
rect 800 140424 453336 142592
rect 880 140144 453336 140424
rect 800 139608 453336 140144
rect 800 139328 453256 139608
rect 800 137976 453336 139328
rect 880 137696 453336 137976
rect 800 135528 453336 137696
rect 880 135248 453336 135528
rect 800 134032 453336 135248
rect 800 133752 453256 134032
rect 800 133080 453336 133752
rect 880 132800 453336 133080
rect 800 130632 453336 132800
rect 880 130352 453336 130632
rect 800 128456 453336 130352
rect 800 128184 453256 128456
rect 880 128176 453256 128184
rect 880 127904 453336 128176
rect 800 125736 453336 127904
rect 880 125456 453336 125736
rect 800 123288 453336 125456
rect 880 123008 453336 123288
rect 800 122880 453336 123008
rect 800 122600 453256 122880
rect 800 120840 453336 122600
rect 880 120560 453336 120840
rect 800 118392 453336 120560
rect 880 118112 453336 118392
rect 800 117304 453336 118112
rect 800 117024 453256 117304
rect 800 115944 453336 117024
rect 880 115664 453336 115944
rect 800 113496 453336 115664
rect 880 113216 453336 113496
rect 800 111728 453336 113216
rect 800 111448 453256 111728
rect 800 111048 453336 111448
rect 880 110768 453336 111048
rect 800 108600 453336 110768
rect 880 108320 453336 108600
rect 800 106152 453336 108320
rect 880 105872 453256 106152
rect 800 103704 453336 105872
rect 880 103424 453336 103704
rect 800 101256 453336 103424
rect 880 100976 453336 101256
rect 800 100576 453336 100976
rect 800 100296 453256 100576
rect 800 98808 453336 100296
rect 880 98528 453336 98808
rect 800 96360 453336 98528
rect 880 96080 453336 96360
rect 800 95000 453336 96080
rect 800 94720 453256 95000
rect 800 93912 453336 94720
rect 880 93632 453336 93912
rect 800 91464 453336 93632
rect 880 91184 453336 91464
rect 800 89424 453336 91184
rect 800 89144 453256 89424
rect 800 89016 453336 89144
rect 880 88736 453336 89016
rect 800 86568 453336 88736
rect 880 86288 453336 86568
rect 800 84120 453336 86288
rect 880 83848 453336 84120
rect 880 83840 453256 83848
rect 800 83568 453256 83840
rect 800 81672 453336 83568
rect 880 81392 453336 81672
rect 800 79224 453336 81392
rect 880 78944 453336 79224
rect 800 78272 453336 78944
rect 800 77992 453256 78272
rect 800 76776 453336 77992
rect 880 76496 453336 76776
rect 800 74328 453336 76496
rect 880 74048 453336 74328
rect 800 72696 453336 74048
rect 800 72416 453256 72696
rect 800 71880 453336 72416
rect 880 71600 453336 71880
rect 800 69432 453336 71600
rect 880 69152 453336 69432
rect 800 67120 453336 69152
rect 800 66984 453256 67120
rect 880 66840 453256 66984
rect 880 66704 453336 66840
rect 800 64536 453336 66704
rect 880 64256 453336 64536
rect 800 62088 453336 64256
rect 880 61808 453336 62088
rect 800 61544 453336 61808
rect 800 61264 453256 61544
rect 800 59640 453336 61264
rect 880 59360 453336 59640
rect 800 57192 453336 59360
rect 880 56912 453336 57192
rect 800 55968 453336 56912
rect 800 55688 453256 55968
rect 800 54744 453336 55688
rect 880 54464 453336 54744
rect 800 52296 453336 54464
rect 880 52016 453336 52296
rect 800 50392 453336 52016
rect 800 50112 453256 50392
rect 800 49848 453336 50112
rect 880 49568 453336 49848
rect 800 47400 453336 49568
rect 880 47120 453336 47400
rect 800 44952 453336 47120
rect 880 44816 453336 44952
rect 880 44672 453256 44816
rect 800 44536 453256 44672
rect 800 42504 453336 44536
rect 880 42224 453336 42504
rect 800 40056 453336 42224
rect 880 39776 453336 40056
rect 800 39240 453336 39776
rect 800 38960 453256 39240
rect 800 37608 453336 38960
rect 880 37328 453336 37608
rect 800 35160 453336 37328
rect 880 34880 453336 35160
rect 800 33664 453336 34880
rect 800 33384 453256 33664
rect 800 32712 453336 33384
rect 880 32432 453336 32712
rect 800 30264 453336 32432
rect 880 29984 453336 30264
rect 800 28088 453336 29984
rect 800 27816 453256 28088
rect 880 27808 453256 27816
rect 880 27536 453336 27808
rect 800 25368 453336 27536
rect 880 25088 453336 25368
rect 800 22920 453336 25088
rect 880 22640 453336 22920
rect 800 22512 453336 22640
rect 800 22232 453256 22512
rect 800 20472 453336 22232
rect 880 20192 453336 20472
rect 800 18024 453336 20192
rect 880 17744 453336 18024
rect 800 16936 453336 17744
rect 800 16656 453256 16936
rect 800 15576 453336 16656
rect 880 15296 453336 15576
rect 800 13128 453336 15296
rect 880 12848 453336 13128
rect 800 11360 453336 12848
rect 800 11080 453256 11360
rect 800 10680 453336 11080
rect 880 10400 453336 10680
rect 800 8232 453336 10400
rect 880 7952 453336 8232
rect 800 5784 453336 7952
rect 800 5504 453256 5784
rect 800 2143 453336 5504
<< metal4 >>
rect 9316 171856 9636 255728
rect 9316 17360 9636 102320
rect 14144 2128 14464 270960
rect 40659 254270 40979 270960
rect 67174 254270 67494 270960
rect 93689 254270 94009 270960
rect 40659 100336 40979 173098
rect 67174 100336 67494 172974
rect 93689 100336 94009 173098
rect 40659 2128 40979 19164
rect 67174 2128 67494 19164
rect 93689 2128 94009 19164
rect 120204 2128 120524 270960
rect 120820 171856 121140 255728
rect 146719 254270 147039 270960
rect 173234 254270 173554 270960
rect 199749 254270 200069 270960
rect 120820 17360 121140 102320
rect 146719 100336 147039 173098
rect 173234 100336 173554 172974
rect 199749 100336 200069 173098
rect 146719 2128 147039 19164
rect 173234 2128 173554 19164
rect 199749 2128 200069 19164
rect 226264 2128 226584 270960
rect 226804 171856 227124 255728
rect 252779 254270 253099 270960
rect 279294 254270 279614 270960
rect 305809 254270 306129 270960
rect 226804 17360 227124 102320
rect 252779 100336 253099 173098
rect 279294 100336 279614 172974
rect 305809 100336 306129 173098
rect 252779 2128 253099 19164
rect 279294 2128 279614 19164
rect 305809 2128 306129 19164
rect 332324 2128 332644 270960
rect 332972 171856 333292 255728
rect 358839 254270 359159 270960
rect 385354 254270 385674 270960
rect 411869 254270 412189 270960
rect 332972 17360 333292 102320
rect 358839 100336 359159 173098
rect 385354 100336 385674 172974
rect 411869 100336 412189 173098
rect 358839 2128 359159 19164
rect 385354 2128 385674 19164
rect 411869 2128 412189 19164
rect 438384 2128 438704 270960
rect 444476 171856 444796 255728
rect 444476 17360 444796 102320
<< obsm4 >>
rect 15699 254190 40579 257141
rect 41059 254190 67094 257141
rect 67574 254190 93609 257141
rect 94089 254190 120124 257141
rect 15699 173178 120124 254190
rect 15699 100256 40579 173178
rect 41059 173054 93609 173178
rect 41059 100256 67094 173054
rect 67574 100256 93609 173054
rect 94089 100256 120124 173178
rect 15699 19244 120124 100256
rect 15699 7923 40579 19244
rect 41059 7923 67094 19244
rect 67574 7923 93609 19244
rect 94089 7923 120124 19244
rect 120604 255808 146639 257141
rect 120604 171776 120740 255808
rect 121220 254190 146639 255808
rect 147119 254190 173154 257141
rect 173634 254190 199669 257141
rect 200149 254190 226184 257141
rect 121220 173178 226184 254190
rect 121220 171776 146639 173178
rect 120604 102400 146639 171776
rect 120604 17280 120740 102400
rect 121220 100256 146639 102400
rect 147119 173054 199669 173178
rect 147119 100256 173154 173054
rect 173634 100256 199669 173054
rect 200149 100256 226184 173178
rect 121220 19244 226184 100256
rect 121220 17280 146639 19244
rect 120604 7923 146639 17280
rect 147119 7923 173154 19244
rect 173634 7923 199669 19244
rect 200149 7923 226184 19244
rect 226664 255808 252699 257141
rect 226664 171776 226724 255808
rect 227204 254190 252699 255808
rect 253179 254190 279214 257141
rect 279694 254190 305729 257141
rect 306209 254190 332244 257141
rect 227204 173178 332244 254190
rect 227204 171776 252699 173178
rect 226664 102400 252699 171776
rect 226664 17280 226724 102400
rect 227204 100256 252699 102400
rect 253179 173054 305729 173178
rect 253179 100256 279214 173054
rect 279694 100256 305729 173054
rect 306209 100256 332244 173178
rect 227204 19244 332244 100256
rect 227204 17280 252699 19244
rect 226664 7923 252699 17280
rect 253179 7923 279214 19244
rect 279694 7923 305729 19244
rect 306209 7923 332244 19244
rect 332724 255808 358759 257141
rect 332724 171776 332892 255808
rect 333372 254190 358759 255808
rect 359239 254190 385274 257141
rect 385754 254190 411789 257141
rect 412269 254190 437493 257141
rect 333372 173178 437493 254190
rect 333372 171776 358759 173178
rect 332724 102400 358759 171776
rect 332724 17280 332892 102400
rect 333372 100256 358759 102400
rect 359239 173054 411789 173178
rect 359239 100256 385274 173054
rect 385754 100256 411789 173054
rect 412269 100256 437493 173178
rect 333372 19244 437493 100256
rect 333372 17280 358759 19244
rect 332724 7923 358759 17280
rect 359239 7923 385274 19244
rect 385754 7923 411789 19244
rect 412269 7923 437493 19244
<< labels >>
rlabel metal4 s 40659 2128 40979 19164 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 40659 100336 40979 173098 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 40659 254270 40979 270960 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 93689 2128 94009 19164 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 93689 100336 94009 173098 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 93689 254270 94009 270960 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 146719 2128 147039 19164 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 146719 100336 147039 173098 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 146719 254270 147039 270960 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 199749 2128 200069 19164 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 199749 100336 200069 173098 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 199749 254270 200069 270960 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252779 2128 253099 19164 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252779 100336 253099 173098 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252779 254270 253099 270960 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 305809 2128 306129 19164 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 305809 100336 306129 173098 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 305809 254270 306129 270960 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 358839 2128 359159 19164 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 358839 100336 359159 173098 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 358839 254270 359159 270960 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 411869 2128 412189 19164 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 411869 100336 412189 173098 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 411869 254270 412189 270960 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 9316 17360 9636 102320 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 120820 171856 121140 255728 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 9316 171856 9636 255728 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 120820 17360 121140 102320 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 226804 17360 227124 102320 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332972 171856 333292 255728 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 226804 171856 227124 255728 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332972 17360 333292 102320 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 444476 17360 444796 102320 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 444476 171856 444796 255728 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 14144 2128 14464 270960 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 67174 2128 67494 19164 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 67174 100336 67494 172974 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 67174 254270 67494 270960 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 120204 2128 120524 270960 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 173234 2128 173554 19164 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 173234 100336 173554 172974 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 173234 254270 173554 270960 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 226264 2128 226584 270960 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 279294 2128 279614 19164 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 279294 100336 279614 172974 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 279294 254270 279614 270960 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 332324 2128 332644 270960 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 385354 2128 385674 19164 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 385354 100336 385674 172974 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 385354 254270 385674 270960 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 438384 2128 438704 270960 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 453336 5584 454136 5704 6 io_in[0]
port 3 nsew signal input
rlabel metal3 s 453336 172864 454136 172984 6 io_in[10]
port 4 nsew signal input
rlabel metal3 s 453336 189592 454136 189712 6 io_in[11]
port 5 nsew signal input
rlabel metal3 s 453336 206320 454136 206440 6 io_in[12]
port 6 nsew signal input
rlabel metal3 s 453336 223048 454136 223168 6 io_in[13]
port 7 nsew signal input
rlabel metal3 s 453336 239776 454136 239896 6 io_in[14]
port 8 nsew signal input
rlabel metal3 s 453336 256504 454136 256624 6 io_in[15]
port 9 nsew signal input
rlabel metal3 s 453336 22312 454136 22432 6 io_in[1]
port 10 nsew signal input
rlabel metal3 s 453336 39040 454136 39160 6 io_in[2]
port 11 nsew signal input
rlabel metal3 s 453336 55768 454136 55888 6 io_in[3]
port 12 nsew signal input
rlabel metal3 s 453336 72496 454136 72616 6 io_in[4]
port 13 nsew signal input
rlabel metal3 s 453336 89224 454136 89344 6 io_in[5]
port 14 nsew signal input
rlabel metal3 s 453336 105952 454136 106072 6 io_in[6]
port 15 nsew signal input
rlabel metal3 s 453336 122680 454136 122800 6 io_in[7]
port 16 nsew signal input
rlabel metal3 s 453336 139408 454136 139528 6 io_in[8]
port 17 nsew signal input
rlabel metal3 s 453336 156136 454136 156256 6 io_in[9]
port 18 nsew signal input
rlabel metal3 s 453336 11160 454136 11280 6 io_oeb[0]
port 19 nsew signal output
rlabel metal3 s 453336 178440 454136 178560 6 io_oeb[10]
port 20 nsew signal output
rlabel metal3 s 453336 195168 454136 195288 6 io_oeb[11]
port 21 nsew signal output
rlabel metal3 s 453336 211896 454136 212016 6 io_oeb[12]
port 22 nsew signal output
rlabel metal3 s 453336 228624 454136 228744 6 io_oeb[13]
port 23 nsew signal output
rlabel metal3 s 453336 245352 454136 245472 6 io_oeb[14]
port 24 nsew signal output
rlabel metal3 s 453336 262080 454136 262200 6 io_oeb[15]
port 25 nsew signal output
rlabel metal3 s 453336 27888 454136 28008 6 io_oeb[1]
port 26 nsew signal output
rlabel metal3 s 453336 44616 454136 44736 6 io_oeb[2]
port 27 nsew signal output
rlabel metal3 s 453336 61344 454136 61464 6 io_oeb[3]
port 28 nsew signal output
rlabel metal3 s 453336 78072 454136 78192 6 io_oeb[4]
port 29 nsew signal output
rlabel metal3 s 453336 94800 454136 94920 6 io_oeb[5]
port 30 nsew signal output
rlabel metal3 s 453336 111528 454136 111648 6 io_oeb[6]
port 31 nsew signal output
rlabel metal3 s 453336 128256 454136 128376 6 io_oeb[7]
port 32 nsew signal output
rlabel metal3 s 453336 144984 454136 145104 6 io_oeb[8]
port 33 nsew signal output
rlabel metal3 s 453336 161712 454136 161832 6 io_oeb[9]
port 34 nsew signal output
rlabel metal3 s 453336 16736 454136 16856 6 io_out[0]
port 35 nsew signal output
rlabel metal3 s 453336 184016 454136 184136 6 io_out[10]
port 36 nsew signal output
rlabel metal3 s 453336 200744 454136 200864 6 io_out[11]
port 37 nsew signal output
rlabel metal3 s 453336 217472 454136 217592 6 io_out[12]
port 38 nsew signal output
rlabel metal3 s 453336 234200 454136 234320 6 io_out[13]
port 39 nsew signal output
rlabel metal3 s 453336 250928 454136 251048 6 io_out[14]
port 40 nsew signal output
rlabel metal3 s 453336 267656 454136 267776 6 io_out[15]
port 41 nsew signal output
rlabel metal3 s 453336 33464 454136 33584 6 io_out[1]
port 42 nsew signal output
rlabel metal3 s 453336 50192 454136 50312 6 io_out[2]
port 43 nsew signal output
rlabel metal3 s 453336 66920 454136 67040 6 io_out[3]
port 44 nsew signal output
rlabel metal3 s 453336 83648 454136 83768 6 io_out[4]
port 45 nsew signal output
rlabel metal3 s 453336 100376 454136 100496 6 io_out[5]
port 46 nsew signal output
rlabel metal3 s 453336 117104 454136 117224 6 io_out[6]
port 47 nsew signal output
rlabel metal3 s 453336 133832 454136 133952 6 io_out[7]
port 48 nsew signal output
rlabel metal3 s 453336 150560 454136 150680 6 io_out[8]
port 49 nsew signal output
rlabel metal3 s 453336 167288 454136 167408 6 io_out[9]
port 50 nsew signal output
rlabel metal2 s 340510 272634 340566 273434 6 one
port 51 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 wb_clk_i
port 52 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 wb_rst_i
port 53 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 wbs_ack_o
port 54 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 wbs_adr_i[0]
port 55 nsew signal input
rlabel metal3 s 0 105952 800 106072 6 wbs_adr_i[10]
port 56 nsew signal input
rlabel metal3 s 0 113296 800 113416 6 wbs_adr_i[11]
port 57 nsew signal input
rlabel metal3 s 0 120640 800 120760 6 wbs_adr_i[12]
port 58 nsew signal input
rlabel metal3 s 0 127984 800 128104 6 wbs_adr_i[13]
port 59 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 wbs_adr_i[14]
port 60 nsew signal input
rlabel metal3 s 0 142672 800 142792 6 wbs_adr_i[15]
port 61 nsew signal input
rlabel metal3 s 0 150016 800 150136 6 wbs_adr_i[16]
port 62 nsew signal input
rlabel metal3 s 0 157360 800 157480 6 wbs_adr_i[17]
port 63 nsew signal input
rlabel metal3 s 0 164704 800 164824 6 wbs_adr_i[18]
port 64 nsew signal input
rlabel metal3 s 0 172048 800 172168 6 wbs_adr_i[19]
port 65 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 wbs_adr_i[1]
port 66 nsew signal input
rlabel metal3 s 0 179392 800 179512 6 wbs_adr_i[20]
port 67 nsew signal input
rlabel metal3 s 0 186736 800 186856 6 wbs_adr_i[21]
port 68 nsew signal input
rlabel metal3 s 0 194080 800 194200 6 wbs_adr_i[22]
port 69 nsew signal input
rlabel metal3 s 0 201424 800 201544 6 wbs_adr_i[23]
port 70 nsew signal input
rlabel metal3 s 0 208768 800 208888 6 wbs_adr_i[24]
port 71 nsew signal input
rlabel metal3 s 0 216112 800 216232 6 wbs_adr_i[25]
port 72 nsew signal input
rlabel metal3 s 0 223456 800 223576 6 wbs_adr_i[26]
port 73 nsew signal input
rlabel metal3 s 0 230800 800 230920 6 wbs_adr_i[27]
port 74 nsew signal input
rlabel metal3 s 0 238144 800 238264 6 wbs_adr_i[28]
port 75 nsew signal input
rlabel metal3 s 0 245488 800 245608 6 wbs_adr_i[29]
port 76 nsew signal input
rlabel metal3 s 0 42304 800 42424 6 wbs_adr_i[2]
port 77 nsew signal input
rlabel metal3 s 0 252832 800 252952 6 wbs_adr_i[30]
port 78 nsew signal input
rlabel metal3 s 0 260176 800 260296 6 wbs_adr_i[31]
port 79 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 wbs_adr_i[3]
port 80 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 wbs_adr_i[4]
port 81 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 wbs_adr_i[5]
port 82 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 wbs_adr_i[6]
port 83 nsew signal input
rlabel metal3 s 0 83920 800 84040 6 wbs_adr_i[7]
port 84 nsew signal input
rlabel metal3 s 0 91264 800 91384 6 wbs_adr_i[8]
port 85 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 wbs_adr_i[9]
port 86 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 wbs_cyc_i
port 87 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 wbs_dat_i[0]
port 88 nsew signal input
rlabel metal3 s 0 108400 800 108520 6 wbs_dat_i[10]
port 89 nsew signal input
rlabel metal3 s 0 115744 800 115864 6 wbs_dat_i[11]
port 90 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 wbs_dat_i[12]
port 91 nsew signal input
rlabel metal3 s 0 130432 800 130552 6 wbs_dat_i[13]
port 92 nsew signal input
rlabel metal3 s 0 137776 800 137896 6 wbs_dat_i[14]
port 93 nsew signal input
rlabel metal3 s 0 145120 800 145240 6 wbs_dat_i[15]
port 94 nsew signal input
rlabel metal3 s 0 152464 800 152584 6 wbs_dat_i[16]
port 95 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 wbs_dat_i[17]
port 96 nsew signal input
rlabel metal3 s 0 167152 800 167272 6 wbs_dat_i[18]
port 97 nsew signal input
rlabel metal3 s 0 174496 800 174616 6 wbs_dat_i[19]
port 98 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 wbs_dat_i[1]
port 99 nsew signal input
rlabel metal3 s 0 181840 800 181960 6 wbs_dat_i[20]
port 100 nsew signal input
rlabel metal3 s 0 189184 800 189304 6 wbs_dat_i[21]
port 101 nsew signal input
rlabel metal3 s 0 196528 800 196648 6 wbs_dat_i[22]
port 102 nsew signal input
rlabel metal3 s 0 203872 800 203992 6 wbs_dat_i[23]
port 103 nsew signal input
rlabel metal3 s 0 211216 800 211336 6 wbs_dat_i[24]
port 104 nsew signal input
rlabel metal3 s 0 218560 800 218680 6 wbs_dat_i[25]
port 105 nsew signal input
rlabel metal3 s 0 225904 800 226024 6 wbs_dat_i[26]
port 106 nsew signal input
rlabel metal3 s 0 233248 800 233368 6 wbs_dat_i[27]
port 107 nsew signal input
rlabel metal3 s 0 240592 800 240712 6 wbs_dat_i[28]
port 108 nsew signal input
rlabel metal3 s 0 247936 800 248056 6 wbs_dat_i[29]
port 109 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 wbs_dat_i[2]
port 110 nsew signal input
rlabel metal3 s 0 255280 800 255400 6 wbs_dat_i[30]
port 111 nsew signal input
rlabel metal3 s 0 262624 800 262744 6 wbs_dat_i[31]
port 112 nsew signal input
rlabel metal3 s 0 54544 800 54664 6 wbs_dat_i[3]
port 113 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 wbs_dat_i[4]
port 114 nsew signal input
rlabel metal3 s 0 71680 800 71800 6 wbs_dat_i[5]
port 115 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 wbs_dat_i[6]
port 116 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 wbs_dat_i[7]
port 117 nsew signal input
rlabel metal3 s 0 93712 800 93832 6 wbs_dat_i[8]
port 118 nsew signal input
rlabel metal3 s 0 101056 800 101176 6 wbs_dat_i[9]
port 119 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 wbs_dat_o[0]
port 120 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 wbs_dat_o[10]
port 121 nsew signal output
rlabel metal3 s 0 118192 800 118312 6 wbs_dat_o[11]
port 122 nsew signal output
rlabel metal3 s 0 125536 800 125656 6 wbs_dat_o[12]
port 123 nsew signal output
rlabel metal3 s 0 132880 800 133000 6 wbs_dat_o[13]
port 124 nsew signal output
rlabel metal3 s 0 140224 800 140344 6 wbs_dat_o[14]
port 125 nsew signal output
rlabel metal3 s 0 147568 800 147688 6 wbs_dat_o[15]
port 126 nsew signal output
rlabel metal3 s 0 154912 800 155032 6 wbs_dat_o[16]
port 127 nsew signal output
rlabel metal3 s 0 162256 800 162376 6 wbs_dat_o[17]
port 128 nsew signal output
rlabel metal3 s 0 169600 800 169720 6 wbs_dat_o[18]
port 129 nsew signal output
rlabel metal3 s 0 176944 800 177064 6 wbs_dat_o[19]
port 130 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 wbs_dat_o[1]
port 131 nsew signal output
rlabel metal3 s 0 184288 800 184408 6 wbs_dat_o[20]
port 132 nsew signal output
rlabel metal3 s 0 191632 800 191752 6 wbs_dat_o[21]
port 133 nsew signal output
rlabel metal3 s 0 198976 800 199096 6 wbs_dat_o[22]
port 134 nsew signal output
rlabel metal3 s 0 206320 800 206440 6 wbs_dat_o[23]
port 135 nsew signal output
rlabel metal3 s 0 213664 800 213784 6 wbs_dat_o[24]
port 136 nsew signal output
rlabel metal3 s 0 221008 800 221128 6 wbs_dat_o[25]
port 137 nsew signal output
rlabel metal3 s 0 228352 800 228472 6 wbs_dat_o[26]
port 138 nsew signal output
rlabel metal3 s 0 235696 800 235816 6 wbs_dat_o[27]
port 139 nsew signal output
rlabel metal3 s 0 243040 800 243160 6 wbs_dat_o[28]
port 140 nsew signal output
rlabel metal3 s 0 250384 800 250504 6 wbs_dat_o[29]
port 141 nsew signal output
rlabel metal3 s 0 47200 800 47320 6 wbs_dat_o[2]
port 142 nsew signal output
rlabel metal3 s 0 257728 800 257848 6 wbs_dat_o[30]
port 143 nsew signal output
rlabel metal3 s 0 265072 800 265192 6 wbs_dat_o[31]
port 144 nsew signal output
rlabel metal3 s 0 56992 800 57112 6 wbs_dat_o[3]
port 145 nsew signal output
rlabel metal3 s 0 66784 800 66904 6 wbs_dat_o[4]
port 146 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 wbs_dat_o[5]
port 147 nsew signal output
rlabel metal3 s 0 81472 800 81592 6 wbs_dat_o[6]
port 148 nsew signal output
rlabel metal3 s 0 88816 800 88936 6 wbs_dat_o[7]
port 149 nsew signal output
rlabel metal3 s 0 96160 800 96280 6 wbs_dat_o[8]
port 150 nsew signal output
rlabel metal3 s 0 103504 800 103624 6 wbs_dat_o[9]
port 151 nsew signal output
rlabel metal3 s 0 30064 800 30184 6 wbs_sel_i[0]
port 152 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 wbs_sel_i[1]
port 153 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 wbs_sel_i[2]
port 154 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 wbs_sel_i[3]
port 155 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 wbs_stb_i
port 156 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 wbs_we_i
port 157 nsew signal input
rlabel metal2 s 113454 272634 113510 273434 6 zero
port 158 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 454136 273434
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 53153936
string GDS_FILE /home/videogamo/Work/mpw8/caravel_pyfive/openlane/pyfive_top/runs/22_12_30_14_40/results/signoff/pyfive_top.magic.gds
string GDS_START 11344096
<< end >>

